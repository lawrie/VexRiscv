`define INCLUDE_QUADRATURE
`define INCLUDE_SEVEN_SEGMENT_A
`define INCLUDE_PULSE_IN
`define INCLUDE_MUX
`define INCLUDE_TONE
`define INCLUDE_SHIFT_OUT
`define INCLUDE_PIN_INTERRUPT
`define INCLUDE_I2C
`define INCLUDE_SHIFT_IN
`define INCLUDE_GPIO_B
`define INCLUDE_UART
`define INCLUDE_SEVEN_SEGMENT_B
`define INCLUDE_SPI_MASTER
`define INCLUDE_WS2811
`define INCLUDE_PS2
`define INCLUDE_QSPI_ANALOG
`define INCLUDE_PWM
`define INCLUDE_GPIO_A
`define INCLUDE_SERVO
`define INCLUDE_TIMER
`define INCLUDE_MACHINE_TIMER

`define MUX_SEVEN_SEGMENT_A 4
`define MUX_TONE 9
`define MUX_SHIFT_OUT 1
`define MUX_SHIFT_IN 0
`define MUX_SEVEN_SEGMENT_B 2
`define MUX_SPI_MASTER 5
`define MUX_WS2811 12
`define MUX_PWM_0  6
`define MUX_PWM_1  7
`define MUX_PWM_2  8
`define MUX_PWM_3  10
`define MUX_PWM_4 11
`define MUX_SERVO 3
