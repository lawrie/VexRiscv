`define GPIO_A_WIDTH 32
`define IO_GPIO_A_WIDTH 32 
`define GPIO_B_WIDTH 17
`define IO_GPIO_B_WIDTH 32 
`define PIN_INTERRUPT_WIDTH 2
`define PWM_WIDTH 5
`define SRAM_ADDRESS_WIDTH 18
`define SRAM_DATA_WIDTH 16

`define INCLUDE_GPIO_A
`define INCLUDE_GPIO_B
`define INCLUDE_I2C
`define INCLUDE_JTAG
`define INCLUDE_MACHINE_TIMER
`define INCLUDE_MUX
`define INCLUDE_PIN_INTERRUPT
`define INCLUDE_PWM
`define INCLUDE_QSPI_ANALOG
`define INCLUDE_SEVEN_SEGMENT_A
`define INCLUDE_SEVEN_SEGMENT_B
`define INCLUDE_SPI_MASTER
`define INCLUDE_SPI_MASTER_A
`define INCLUDE_SRAM
`define INCLUDE_TIMER
`define INCLUDE_UART
`define INCLUDE_UART_A
`define INCLUDE_WS2811

`define MUX_PWM_0 6
`define MUX_PWM_1 7
`define MUX_PWM_2 8
`define MUX_PWM_3 10
`define MUX_PWM_4 11
`define MUX_SEVEN_SEGMENT_A 4
`define MUX_SEVEN_SEGMENT_B 2
`define MUX_SPI_MASTER 5
`define MUX_SPI_MASTER_A 14
`define MUX_UART_A 13
`define MUX_WS2811 12
